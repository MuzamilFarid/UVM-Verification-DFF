
class dff-test extends uvm_test;





endclass